`default_nettype none

module \std::cdc::sync2_bool  (
        input clk_i,
        input in_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::cdc::sync2_bool" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::cdc::sync2_bool );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/cdc.spade:34,9" *)
    logic _e_136;
    (* src = "<compiler dir>/stdlib/cdc.spade:34,9" *)
    \std::cdc::sync2[565]  sync2_0(.clk_i(\clk ), .in_i(\in ), .output__(_e_136));
    assign output__ = _e_136;
endmodule

module \std::conv::bit_to_bool  (
        input b_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::bit_to_bool" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::bit_to_bool );
        end
    end
    `endif
    logic \b ;
    assign \b  = b_i;
    logic _e_432;
    assign _e_432 = \b ;
    assign output__ = _e_432;
endmodule

module \std::conv::clock_to_bool  (
        input c_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::clock_to_bool" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::clock_to_bool );
        end
    end
    `endif
    logic \c ;
    assign \c  = c_i;
    logic _e_486;
    assign _e_486 = \c ;
    assign output__ = _e_486;
endmodule

module \std::conv::bool_to_clock  (
        input c_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::bool_to_clock" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::bool_to_clock );
        end
    end
    `endif
    logic \c ;
    assign \c  = c_i;
    logic _e_490;
    assign _e_490 = \c ;
    assign output__ = _e_490;
endmodule

module \std::io::rising_edge  (
        input clk_i,
        input sync1_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::io::rising_edge" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::io::rising_edge );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \sync1 ;
    assign \sync1  = sync1_i;
    (* src = "<compiler dir>/stdlib/io.spade:3,14" *)
    reg \sync2 ;
    (* src = "<compiler dir>/stdlib/io.spade:4,14" *)
    logic _e_574;
    (* src = "<compiler dir>/stdlib/io.spade:4,5" *)
    logic _e_572;
    always @(posedge \clk ) begin
        \sync2  <= \sync1 ;
    end
    assign _e_574 = !\sync2 ;
    assign _e_572 = \sync1  && _e_574;
    assign output__ = _e_572;
endmodule

module \std::io::falling_edge  (
        input clk_i,
        input sync1_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::io::falling_edge" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::io::falling_edge );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \sync1 ;
    assign \sync1  = sync1_i;
    (* src = "<compiler dir>/stdlib/io.spade:9,14" *)
    reg \sync2 ;
    (* src = "<compiler dir>/stdlib/io.spade:10,14" *)
    logic _e_582;
    (* src = "<compiler dir>/stdlib/io.spade:10,5" *)
    logic _e_580;
    always @(posedge \clk ) begin
        \sync2  <= \sync1 ;
    end
    assign _e_582 = !\sync1 ;
    assign _e_580 = \sync2  && _e_582;
    assign output__ = _e_580;
endmodule

module \swim_tinytapeout::design  (
        input clk_i,
        input rst_i,
        input[7:0] ui_in_i,
        output[7:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "swim_tinytapeout::design" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \swim_tinytapeout::design );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \rst ;
    assign \rst  = rst_i;
    logic[7:0] \ui_in ;
    assign \ui_in  = ui_in_i;
    (* src = "src/main.spade:4,58" *)
    logic _e_1082;
    (* src = "src/main.spade:7,15" *)
    logic[32:0] _e_1089;
    (* src = "src/main.spade:7,9" *)
    logic[31:0] _e_1088;
    (* src = "src/main.spade:4,55" *)
    logic[31:0] _e_1081;
    (* src = "src/main.spade:4,14" *)
    reg[31:0] \second_counter ;
    (* src = "src/main.spade:11,37" *)
    logic _e_1097;
    (* src = "src/main.spade:13,13" *)
    logic _e_1103;
    (* src = "src/main.spade:13,12" *)
    logic _e_1102;
    (* src = "src/main.spade:14,19" *)
    logic[8:0] _e_1108;
    (* src = "src/main.spade:14,13" *)
    logic[7:0] _e_1107;
    (* src = "src/main.spade:16,19" *)
    logic[8:0] _e_1113;
    (* src = "src/main.spade:16,13" *)
    logic[7:0] _e_1112;
    (* src = "src/main.spade:13,9" *)
    logic[7:0] _e_1101;
    (* src = "src/main.spade:11,34" *)
    logic[7:0] _e_1096;
    (* src = "src/main.spade:11,14" *)
    reg[7:0] \val ;
    localparam[31:0] _e_1080 = 32'd0;
    localparam[31:0] _e_1084 = 32'd1000;
    assign _e_1082 = \second_counter  == _e_1084;
    localparam[31:0] _e_1086 = 32'd0;
    localparam[31:0] _e_1091 = 32'd1;
    assign _e_1089 = \second_counter  + _e_1091;
    assign _e_1088 = _e_1089[31:0];
    assign _e_1081 = _e_1082 ? _e_1086 : _e_1088;
    always @(posedge \clk ) begin
        if (\rst ) begin
            \second_counter  <= _e_1080;
        end
        else begin
            \second_counter  <= _e_1081;
        end
    end
    localparam[7:0] _e_1095 = 0;
    localparam[31:0] _e_1099 = 32'd0;
    assign _e_1097 = \second_counter  == _e_1099;
    localparam[2:0] _e_1105 = 0;
    assign _e_1103 = \ui_in [_e_1105];
    assign _e_1102 = !_e_1103;
    localparam[7:0] _e_1110 = 1;
    assign _e_1108 = \val  + _e_1110;
    assign _e_1107 = _e_1108[7:0];
    localparam[7:0] _e_1115 = 1;
    assign _e_1113 = \val  - _e_1115;
    assign _e_1112 = _e_1113[7:0];
    assign _e_1101 = _e_1102 ? _e_1107 : _e_1112;
    assign _e_1096 = _e_1097 ? _e_1101 : \val ;
    always @(posedge \clk ) begin
        if (\rst ) begin
            \val  <= _e_1095;
        end
        else begin
            \val  <= _e_1096;
        end
    end
    assign output__ = \val ;
endmodule

module tt_um_your_design (
        input clk,
        input rst_n,
        input[7:0] ui_in,
        output[7:0] uo_out,
        input[7:0] uio_in,
        output[7:0] uio_out,
        output[7:0] uio_oe,
        input ena
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tt_um_your_design" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, tt_um_your_design);
        end
    end
    `endif
    logic[7:0] \uo_out_mut ;
    assign uo_out = \uo_out_mut ;
    logic[7:0] \uio_out_mut ;
    assign uio_out = \uio_out_mut ;
    logic[7:0] \uio_oe_mut ;
    assign uio_oe = \uio_oe_mut ;
    (* src = "src/main.spade:42,15" *)
    logic \rst ;
    (* src = "src/main.spade:44,19" *)
    logic[7:0] _e_1124;
    (* src = "src/main.spade:45,18" *)
    logic[7:0] _e_1127;
    (* src = "src/main.spade:49,18" *)
    logic[7:0] \output ;
    (* src = "src/main.spade:51,19" *)
    logic[7:0] _e_1135;
    assign \rst  = !\rst_n ;
    localparam[7:0] _e_1125 = 0;
    assign _e_1124 = _e_1125;
    assign \uio_out_mut  = _e_1124;
    localparam[7:0] _e_1128 = 0;
    assign _e_1127 = _e_1128;
    assign \uio_oe_mut  = _e_1127;
    (* src = "src/main.spade:49,18" *)
    \swim_tinytapeout::design  design_0(.clk_i(\clk ), .rst_i(\rst ), .ui_in_i(\ui_in ), .output__(\output ));
    (* src = "src/main.spade:51,19" *)
    \std::conv::impl_3::to_bits[566]  to_bits_0(.self_i(\output ), .output__(_e_1135));
    assign \uo_out_mut  = _e_1135;
endmodule

module top (
        input clk,
        input rst_n,
        input[7:0] ui_in,
        output[7:0] uo_out,
        input[7:0] uio_in,
        output[7:0] uio_out,
        output[7:0] uio_oe,
        input ena
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "top" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, top);
        end
    end
    `endif
    logic[7:0] \uo_out_mut ;
    assign uo_out = \uo_out_mut ;
    logic[7:0] \uio_out_mut ;
    assign uio_out = \uio_out_mut ;
    logic[7:0] \uio_oe_mut ;
    assign uio_oe = \uio_oe_mut ;
    (* src = "src/main.spade:68,5" *)
    tt_um_your_design tt_um_your_design_0(.clk(\clk ), .rst_n(\rst_n ), .ui_in(\ui_in ), .uo_out(\uo_out_mut ), .uio_in(\uio_in ), .uio_out(\uio_out_mut ), .uio_oe(\uio_oe_mut ), .ena(\ena ));
endmodule

module \std::conv::impl_4::to_be_bytes  (
        input[15:0] self_i,
        output[15:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::impl_4::to_be_bytes" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::impl_4::to_be_bytes );
        end
    end
    `endif
    logic[15:0] \self ;
    assign \self  = self_i;
    (* src = "<compiler dir>/stdlib/conv.spade:169,16" *)
    logic[15:0] _e_513;
    (* src = "<compiler dir>/stdlib/conv.spade:169,10" *)
    logic[7:0] _e_512;
    (* src = "<compiler dir>/stdlib/conv.spade:169,28" *)
    logic[7:0] _e_516;
    (* src = "<compiler dir>/stdlib/conv.spade:169,9" *)
    logic[15:0] _e_511;
    localparam[15:0] _e_515 = 8;
    assign _e_513 = \self  >> _e_515;
    assign _e_512 = _e_513[7:0];
    assign _e_516 = \self [7:0];
    assign _e_511 = {_e_516, _e_512};
    assign output__ = _e_511;
endmodule

module \std::conv::impl_4::to_le_bytes  (
        input[15:0] self_i,
        output[15:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::impl_4::to_le_bytes" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::impl_4::to_le_bytes );
        end
    end
    `endif
    logic[15:0] \self ;
    assign \self  = self_i;
    (* src = "<compiler dir>/stdlib/conv.spade:175,31" *)
    logic[15:0] _e_520;
    (* src = "<compiler dir>/stdlib/conv.spade:175,9" *)
    logic[15:0] _e_519;
    (* src = "<compiler dir>/stdlib/conv.spade:175,31" *)
    \std::conv::impl_4::to_be_bytes  to_be_bytes_0(.self_i(\self ), .output__(_e_520));
    (* src = "<compiler dir>/stdlib/conv.spade:175,9" *)
    \std::conv::flip_array[567]  flip_array_0(.in_i(_e_520), .output__(_e_519));
    assign output__ = _e_519;
endmodule

module \std::conv::impl_5::to_be_bytes  (
        input[23:0] self_i,
        output[23:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::impl_5::to_be_bytes" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::impl_5::to_be_bytes );
        end
    end
    `endif
    logic[23:0] \self ;
    assign \self  = self_i;
    (* src = "<compiler dir>/stdlib/conv.spade:183,16" *)
    logic[23:0] _e_525;
    (* src = "<compiler dir>/stdlib/conv.spade:183,10" *)
    logic[7:0] _e_524;
    (* src = "<compiler dir>/stdlib/conv.spade:183,35" *)
    logic[23:0] _e_529;
    (* src = "<compiler dir>/stdlib/conv.spade:183,29" *)
    logic[7:0] _e_528;
    (* src = "<compiler dir>/stdlib/conv.spade:183,47" *)
    logic[7:0] _e_532;
    (* src = "<compiler dir>/stdlib/conv.spade:183,9" *)
    logic[23:0] _e_523;
    localparam[23:0] _e_527 = 16;
    assign _e_525 = \self  >> _e_527;
    assign _e_524 = _e_525[7:0];
    localparam[23:0] _e_531 = 8;
    assign _e_529 = \self  >> _e_531;
    assign _e_528 = _e_529[7:0];
    assign _e_532 = \self [7:0];
    assign _e_523 = {_e_532, _e_528, _e_524};
    assign output__ = _e_523;
endmodule

module \std::conv::impl_5::to_le_bytes  (
        input[23:0] self_i,
        output[23:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::impl_5::to_le_bytes" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::impl_5::to_le_bytes );
        end
    end
    `endif
    logic[23:0] \self ;
    assign \self  = self_i;
    (* src = "<compiler dir>/stdlib/conv.spade:189,31" *)
    logic[23:0] _e_536;
    (* src = "<compiler dir>/stdlib/conv.spade:189,9" *)
    logic[23:0] _e_535;
    (* src = "<compiler dir>/stdlib/conv.spade:189,31" *)
    \std::conv::impl_5::to_be_bytes  to_be_bytes_0(.self_i(\self ), .output__(_e_536));
    (* src = "<compiler dir>/stdlib/conv.spade:189,9" *)
    \std::conv::flip_array[568]  flip_array_0(.in_i(_e_536), .output__(_e_535));
    assign output__ = _e_535;
endmodule

module \std::conv::impl_6::to_be_bytes  (
        input[31:0] self_i,
        output[31:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::impl_6::to_be_bytes" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::impl_6::to_be_bytes );
        end
    end
    `endif
    logic[31:0] \self ;
    assign \self  = self_i;
    (* src = "<compiler dir>/stdlib/conv.spade:197,16" *)
    logic[31:0] _e_541;
    (* src = "<compiler dir>/stdlib/conv.spade:197,10" *)
    logic[7:0] _e_540;
    (* src = "<compiler dir>/stdlib/conv.spade:197,35" *)
    logic[31:0] _e_545;
    (* src = "<compiler dir>/stdlib/conv.spade:197,29" *)
    logic[7:0] _e_544;
    (* src = "<compiler dir>/stdlib/conv.spade:197,54" *)
    logic[31:0] _e_549;
    (* src = "<compiler dir>/stdlib/conv.spade:197,48" *)
    logic[7:0] _e_548;
    (* src = "<compiler dir>/stdlib/conv.spade:197,66" *)
    logic[7:0] _e_552;
    (* src = "<compiler dir>/stdlib/conv.spade:197,9" *)
    logic[31:0] _e_539;
    localparam[31:0] _e_543 = 32'd24;
    assign _e_541 = \self  >> _e_543;
    assign _e_540 = _e_541[7:0];
    localparam[31:0] _e_547 = 32'd16;
    assign _e_545 = \self  >> _e_547;
    assign _e_544 = _e_545[7:0];
    localparam[31:0] _e_551 = 32'd8;
    assign _e_549 = \self  >> _e_551;
    assign _e_548 = _e_549[7:0];
    assign _e_552 = \self [7:0];
    assign _e_539 = {_e_552, _e_548, _e_544, _e_540};
    assign output__ = _e_539;
endmodule

module \std::conv::impl_6::to_le_bytes  (
        input[31:0] self_i,
        output[31:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::impl_6::to_le_bytes" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::impl_6::to_le_bytes );
        end
    end
    `endif
    logic[31:0] \self ;
    assign \self  = self_i;
    (* src = "<compiler dir>/stdlib/conv.spade:203,31" *)
    logic[31:0] _e_556;
    (* src = "<compiler dir>/stdlib/conv.spade:203,9" *)
    logic[31:0] _e_555;
    (* src = "<compiler dir>/stdlib/conv.spade:203,31" *)
    \std::conv::impl_6::to_be_bytes  to_be_bytes_0(.self_i(\self ), .output__(_e_556));
    (* src = "<compiler dir>/stdlib/conv.spade:203,9" *)
    \std::conv::flip_array[569]  flip_array_0(.in_i(_e_556), .output__(_e_555));
    assign output__ = _e_555;
endmodule

module \std::cdc::sync2[565]  (
        input clk_i,
        input in_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::cdc::sync2[565]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::cdc::sync2[565] );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/cdc.spade:16,14" *)
    reg \sync1 ;
    (* src = "<compiler dir>/stdlib/cdc.spade:17,14" *)
    reg \sync2 ;
    always @(posedge \clk ) begin
        \sync1  <= \in ;
    end
    always @(posedge \clk ) begin
        \sync2  <= \sync1 ;
    end
    assign output__ = \sync2 ;
endmodule

module \std::conv::impl_3::to_bits[566]  (
        input[7:0] self_i,
        output[7:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::impl_3::to_bits[566]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::impl_3::to_bits[566] );
        end
    end
    `endif
    logic[7:0] \self ;
    assign \self  = self_i;
    (* src = "<compiler dir>/stdlib/conv.spade:160,9" *)
    logic[7:0] _e_508;
    (* src = "<compiler dir>/stdlib/conv.spade:160,9" *)
    \std::conv::uint_to_bits[570]  uint_to_bits_0(.input_i(\self ), .output__(_e_508));
    assign output__ = _e_508;
endmodule

module \std::conv::flip_array[567]  (
        input[15:0] in_i,
        output[15:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::flip_array[567]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::flip_array[567] );
        end
    end
    `endif
    logic[15:0] \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/conv.spade:39,49" *)
    logic[15:0] \result ;
    (* src = "<compiler dir>/stdlib/conv.spade:39,49" *)
    \std::conv::std::conv::flip_array::F[571]  F_0(.in_i(\in ), .output__(\result ));
    assign output__ = \result ;
endmodule

module \std::conv::flip_array[568]  (
        input[23:0] in_i,
        output[23:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::flip_array[568]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::flip_array[568] );
        end
    end
    `endif
    logic[23:0] \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/conv.spade:39,49" *)
    logic[23:0] \result ;
    (* src = "<compiler dir>/stdlib/conv.spade:39,49" *)
    \std::conv::std::conv::flip_array::F[572]  F_0(.in_i(\in ), .output__(\result ));
    assign output__ = \result ;
endmodule

module \std::conv::flip_array[569]  (
        input[31:0] in_i,
        output[31:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::flip_array[569]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::flip_array[569] );
        end
    end
    `endif
    logic[31:0] \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/conv.spade:39,49" *)
    logic[31:0] \result ;
    (* src = "<compiler dir>/stdlib/conv.spade:39,49" *)
    \std::conv::std::conv::flip_array::F[573]  F_0(.in_i(\in ), .output__(\result ));
    assign output__ = \result ;
endmodule

module \std::conv::uint_to_bits[570]  (
        input[7:0] input_i,
        output[7:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::uint_to_bits[570]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::uint_to_bits[570] );
        end
    end
    `endif
    logic[7:0] \input ;
    assign \input  = input_i;
    logic[7:0] _e_470;
    assign _e_470 = \input ;
    assign output__ = _e_470;
endmodule

module \std::conv::std::conv::flip_array::F[571]  (
        input[15:0] in_i,
        output[15:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::std::conv::flip_array::F[571]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::std::conv::flip_array::F[571] );
        end
    end
    `endif
    logic[15:0] \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/conv.spade:43,9" *)
    logic[7:0] _e_440;
    (* src = "<compiler dir>/stdlib/conv.spade:43,47" *)
    logic[7:0] _e_445;
    (* src = "<compiler dir>/stdlib/conv.spade:43,36" *)
    logic[7:0] _e_444;
    (* src = "<compiler dir>/stdlib/conv.spade:43,9" *)
    logic[15:0] _e_439;
    assign _e_440 = \in [15-:8];
    assign _e_445 = \in [7-:8];
    (* src = "<compiler dir>/stdlib/conv.spade:43,36" *)
    \std::conv::flip_array[574]  flip_array_0(.in_i(_e_445), .output__(_e_444));
    (* src = "<compiler dir>/stdlib/conv.spade:43,9" *)
    \std::conv::concat_arrays[575]  concat_arrays_0(.l_i(_e_440), .r_i(_e_444), .output__(_e_439));
    assign output__ = _e_439;
endmodule

module \std::conv::std::conv::flip_array::F[572]  (
        input[23:0] in_i,
        output[23:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::std::conv::flip_array::F[572]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::std::conv::flip_array::F[572] );
        end
    end
    `endif
    logic[23:0] \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/conv.spade:43,9" *)
    logic[7:0] _e_440;
    (* src = "<compiler dir>/stdlib/conv.spade:43,47" *)
    logic[15:0] _e_445;
    (* src = "<compiler dir>/stdlib/conv.spade:43,36" *)
    logic[15:0] _e_444;
    (* src = "<compiler dir>/stdlib/conv.spade:43,9" *)
    logic[23:0] _e_439;
    assign _e_440 = \in [23-:8];
    assign _e_445 = \in [15-:16];
    (* src = "<compiler dir>/stdlib/conv.spade:43,36" *)
    \std::conv::flip_array[567]  flip_array_0(.in_i(_e_445), .output__(_e_444));
    (* src = "<compiler dir>/stdlib/conv.spade:43,9" *)
    \std::conv::concat_arrays[576]  concat_arrays_0(.l_i(_e_440), .r_i(_e_444), .output__(_e_439));
    assign output__ = _e_439;
endmodule

module \std::conv::std::conv::flip_array::F[573]  (
        input[31:0] in_i,
        output[31:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::std::conv::flip_array::F[573]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::std::conv::flip_array::F[573] );
        end
    end
    `endif
    logic[31:0] \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/conv.spade:43,9" *)
    logic[7:0] _e_440;
    (* src = "<compiler dir>/stdlib/conv.spade:43,47" *)
    logic[23:0] _e_445;
    (* src = "<compiler dir>/stdlib/conv.spade:43,36" *)
    logic[23:0] _e_444;
    (* src = "<compiler dir>/stdlib/conv.spade:43,9" *)
    logic[31:0] _e_439;
    assign _e_440 = \in [31-:8];
    assign _e_445 = \in [23-:24];
    (* src = "<compiler dir>/stdlib/conv.spade:43,36" *)
    \std::conv::flip_array[568]  flip_array_0(.in_i(_e_445), .output__(_e_444));
    (* src = "<compiler dir>/stdlib/conv.spade:43,9" *)
    \std::conv::concat_arrays[577]  concat_arrays_0(.l_i(_e_440), .r_i(_e_444), .output__(_e_439));
    assign output__ = _e_439;
endmodule

module \std::conv::flip_array[574]  (
        input[7:0] in_i,
        output[7:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::flip_array[574]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::flip_array[574] );
        end
    end
    `endif
    logic[7:0] \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/conv.spade:39,49" *)
    logic[7:0] \result ;
    (* src = "<compiler dir>/stdlib/conv.spade:39,49" *)
    \std::conv::std::conv::flip_array::F[578]  F_0(.in_i(\in ), .output__(\result ));
    assign output__ = \result ;
endmodule

module \std::conv::concat_arrays[575]  (
        input[7:0] l_i,
        input[7:0] r_i,
        output[15:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::concat_arrays[575]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::concat_arrays[575] );
        end
    end
    `endif
    logic[7:0] \l ;
    assign \l  = l_i;
    logic[7:0] \r ;
    assign \r  = r_i;
    (* src = "<compiler dir>/stdlib/conv.spade:25,30" *)
    logic[15:0] _e_427;
    logic[15:0] _e_426;
    assign _e_427 = {\r , \l };
    assign _e_426 = _e_427;
    assign output__ = _e_426;
endmodule

module \std::conv::concat_arrays[576]  (
        input[7:0] l_i,
        input[15:0] r_i,
        output[23:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::concat_arrays[576]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::concat_arrays[576] );
        end
    end
    `endif
    logic[7:0] \l ;
    assign \l  = l_i;
    logic[15:0] \r ;
    assign \r  = r_i;
    (* src = "<compiler dir>/stdlib/conv.spade:25,30" *)
    logic[23:0] _e_427;
    logic[23:0] _e_426;
    assign _e_427 = {\r , \l };
    assign _e_426 = _e_427;
    assign output__ = _e_426;
endmodule

module \std::conv::concat_arrays[577]  (
        input[7:0] l_i,
        input[23:0] r_i,
        output[31:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::concat_arrays[577]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::concat_arrays[577] );
        end
    end
    `endif
    logic[7:0] \l ;
    assign \l  = l_i;
    logic[23:0] \r ;
    assign \r  = r_i;
    (* src = "<compiler dir>/stdlib/conv.spade:25,30" *)
    logic[31:0] _e_427;
    logic[31:0] _e_426;
    assign _e_427 = {\r , \l };
    assign _e_426 = _e_427;
    assign output__ = _e_426;
endmodule

module \std::conv::std::conv::flip_array::F[578]  (
        input[7:0] in_i,
        output[7:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::std::conv::flip_array::F[578]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::std::conv::flip_array::F[578] );
        end
    end
    `endif
    logic[7:0] \in ;
    assign \in  = in_i;
    (* src = "<compiler dir>/stdlib/conv.spade:43,9" *)
    logic[7:0] _e_440;
    (* src = "<compiler dir>/stdlib/conv.spade:43,9" *)
    logic[7:0] _e_439;
    assign _e_440 = \in ;
    
    (* src = "<compiler dir>/stdlib/conv.spade:43,36" *)
    \std::conv::flip_array[579]  flip_array_0();
    (* src = "<compiler dir>/stdlib/conv.spade:43,9" *)
    \std::conv::concat_arrays[580]  concat_arrays_0(.l_i(_e_440), .output__(_e_439));
    assign output__ = _e_439;
endmodule

module \std::conv::flip_array[579]  (
        
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::flip_array[579]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::flip_array[579] );
        end
    end
    `endif
    (* src = "<compiler dir>/stdlib/conv.spade:39,49" *)
    \std::conv::std::conv::flip_array::T[581]  T_0();
endmodule

module \std::conv::concat_arrays[580]  (
        input[7:0] l_i,
        output[7:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::concat_arrays[580]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::concat_arrays[580] );
        end
    end
    `endif
    logic[7:0] \l ;
    assign \l  = l_i;
    (* src = "<compiler dir>/stdlib/conv.spade:25,30" *)
    logic[7:0] _e_427;
    logic[7:0] _e_426;
    assign _e_427 = {\l };
    assign _e_426 = _e_427;
    assign output__ = _e_426;
endmodule

module \std::conv::std::conv::flip_array::T[581]  (
        
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::conv::std::conv::flip_array::T[581]" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::conv::std::conv::flip_array::T[581] );
        end
    end
    `endif
    
endmodule